`include "mycpu.h"

module id_stage(
    input                          clk           ,
    input                          reset         ,
    //allowin
    input                          es_allowin    ,
    output                         ds_allowin    ,
    //from fs
    input                          fs_to_ds_valid,
    input  [`FS_TO_DS_BUS_WD -1:0] fs_to_ds_bus  ,
    //to es
    output                         ds_to_es_valid,
    output [`DS_TO_ES_BUS_WD -1:0] ds_to_es_bus  ,
    //to fs
    output [`BR_BUS_WD       -1:0] br_bus        ,
    //to rf: for write back
    input  [`WS_TO_RF_BUS_WD -1:0] ws_to_rf_bus  ,
    //forward valid signal and dest
    input  [`ES_DEST_BUS     -1:0] es_dest_bus   ,
    input  [`MS_DEST_BUS     -1:0] ms_dest_bus   ,
    input  [`WS_DEST_BUS     -1:0] ws_dest_bus   ,
    //forward data
    input  [`ES_TO_DS_BUS    -1:0] es_to_ds_bus  ,
    input  [`MS_TO_DS_BUS    -1:0] ms_to_ds_bus  ,
    input  [`WS_TO_DS_BUS    -1:0] ws_to_ds_bus  ,
    //flush
    input                         ws_flush_ds_bus,
    //interrupt
    input                         has_int
);

reg         ds_valid   ;
wire        ds_ready_go;

reg  [`FS_TO_DS_BUS_WD -1:0] fs_to_ds_bus_r;

wire [31:0] ds_inst;
wire [31:0] ds_pc  ;

wire        ex_ADEF;
wire        ex_INE;
wire        tlb_refill;
wire        inst_page_fault;
wire        plv_illegal;
wire        fs_mmu_ex;

assign {fs_mmu_ex,
        tlb_refill,
        inst_page_fault,
        plv_illegal,
        ex_ADEF,
        ds_inst,
        ds_pc  } = fs_to_ds_bus_r;

wire        rf_we   ;
wire [ 4:0] rf_waddr;
wire [31:0] rf_wdata;
assign {rf_we   ,  //37:37
        rf_waddr,  //36:32
        rf_wdata   //31:0
       } = ws_to_rf_bus;

wire        br_inst_valid;
wire        br_stall;
wire        br_taken;
wire [31:0] br_target;

wire [18:0] alu_op;
wire        src1_is_pc;
wire        src2_is_imm;
wire        res_from_mem;
wire        dst_is_r1;
wire        gr_we;
wire        mem_we;
wire        src_reg_is_rd;
wire [4: 0] dest;
wire [31:0] rj_value;
wire [31:0] rkd_value;
wire [31:0] ds_imm;
wire [31:0] br_offs;
wire [31:0] jirl_offs;

wire rj_le_rd;

wire [ 5:0] op_31_26;
wire [ 3:0] op_25_22;
wire [ 1:0] op_21_20;
wire [ 4:0] op_19_15;
wire [ 4:0] rd;
wire [ 4:0] rj;
wire [ 4:0] rk;
wire [11:0] i12;
wire [19:0] i20;
wire [15:0] i16;
wire [25:0] i26;

wire [63:0] op_31_26_d;
wire [15:0] op_25_22_d;
wire [ 3:0] op_21_20_d;
wire [31:0] op_19_15_d;
  
wire        inst_add_w; 
wire        inst_sub_w;  
wire        inst_slt;    
wire        inst_sltu; 
wire        inst_slti;
wire        inst_sltui;  
wire        inst_nor;    
wire        inst_and;    
wire        inst_or;     
wire        inst_xor; 
wire        inst_andi;
wire        inst_ori;
wire        inst_xori;   
wire        inst_slli_w;  
wire        inst_srli_w;  
wire        inst_srai_w; 
wire        inst_sll_w;
wire        inst_srl_w;
wire        inst_sra_w; 
wire        inst_addi_w; 
wire        inst_ld_w; 
wire        inst_ld_b;
wire        inst_ld_h;
wire        inst_ld_bu;
wire        inst_ld_hu; 
wire        inst_st_w;
wire        inst_st_b;
wire        inst_st_h;   
wire        inst_jirl;   
wire        inst_b;      
wire        inst_bl;     
wire        inst_beq;    
wire        inst_bne;
wire        inst_blt;
wire        inst_bge;
wire        inst_bltu;
wire        inst_bgeu;    
wire        inst_lu12i_w;
wire        inst_pcaddu12i;
wire        inst_mul_w;
wire        inst_mulh_w;
wire        inst_mulh_wu;
wire        inst_div_w;
wire        inst_mod_w;
wire        inst_div_wu;
wire        inst_mod_wu;

//kernel inst
wire        inst_csrrd;
wire        inst_csrwr;
wire        inst_csrxchg;
wire        inst_ertn;
wire        inst_syscall;
wire        inst_break;
wire        inst_rdcntid_w;
wire        inst_rdcntvl_w;
wire        inst_rdcntvh_w;

wire        inst_tlbsrch;
wire        inst_tlbrd;
wire        inst_tlbwr;
wire        inst_tlbfill;
wire        inst_invtlb;

wire        need_ui5;
wire        need_ui12;
wire        need_si12;
wire        need_si16;
wire        need_si20;
wire        need_si26;  
wire        src2_is_4;

wire [ 4:0] rf_raddr1;
wire [31:0] rf_rdata1;
wire [ 4:0] rf_raddr2;
wire [31:0] rf_rdata2;

wire        es_inst_load;
wire        raddr1_valid;
wire        raddr2_valid;
wire        es_read_except;
wire        es_dest_valid;
wire        ms_read_except;
wire        ms_dest_valid;
wire        ws_dest_valid;
wire [ 4:0] es_dest;
wire [ 4:0] ms_dest;
wire [ 4:0] ws_dest;

wire        es_relate_r1;
wire        es_relate_r2;
wire        ms_relate_r1;
wire        ms_relate_r2;
wire        ws_relate_r1;
wire        ws_relate_r2;

wire        es_read1_unuse;
wire        es_read2_unuse;
wire        ms_read1_unuse;
wire        ms_read2_unuse;
wire [ 2:0] inst_st_op;
wire [ 4:0] inst_ld_op;
wire [ 2:0] inst_cnt_op;

wire csr_we;
wire csr_re;
wire [31:0]csr_wmask;
wire [13:0]csr_num;//csr regs number:csrrd csrwr csrxchg
//assign csr_num = inst_ertn ? `CSR_ERA:ds_inst[23:10];//ertn : csr_era

assign {es_inst_load,
        es_read_except,
        es_dest_valid,
        es_dest
       } = es_dest_bus;

assign {ms_read_except,
        ms_dest_valid,
        ms_dest
       } = ms_dest_bus;

assign {ws_dest_valid,
        ws_dest
       } = ws_dest_bus;

wire        rj_eq_rd;
wire        rj_leu_rd;
wire   [4:0]invtlb_op;
wire   [4:0]tlbop;
assign br_bus       = {br_stall,br_taken,br_target};

assign ds_to_es_bus = {fs_mmu_ex,     //235:235
                       tlb_refill,    //234:234
                       inst_page_fault,//233:233
                       plv_illegal,   //232:232
                       tlbop       ,  //231:227  
                       invtlb_op   ,  //226:222
                       inst_cnt_op ,  //221:219
                       has_int     ,  //218:218
                       ex_INE      ,  //217:217
                       ex_ADEF     ,  //216:216
                       inst_break  ,  //215:215
                       inst_ertn   ,  //214:214
                       inst_syscall,  //213:213
                       csr_we      ,  //212:212
                       csr_re      ,  //211:211 
                       csr_wmask   ,  //210:179
                       csr_num     ,  //178:165
                       inst_st_op  ,  //164:162
                       inst_ld_op  ,  //161:157
                       alu_op      ,  //156:138
                       res_from_mem,  //137:137
                       src1_is_pc  ,  //136:136
                       src2_is_imm ,  //135:135
                       gr_we       ,  //134:134
                       mem_we      ,  //133:133
                       dest        ,  //132:128
                       ds_imm      ,  //127:96
                       rj_value    ,  //95 :64
                       rkd_value   ,  //63 :32
                       ds_pc          //31 :0
                      };


assign ds_allowin     = !ds_valid || ds_ready_go && es_allowin;
assign ds_to_es_valid = ds_valid && ds_ready_go;// && !ws_flush_ds_bus;
always @(posedge clk) begin
    if (reset) begin
        ds_valid <= 1'b0;
    end
    else if (/*(br_taken & es_allowin)*/ ws_flush_ds_bus ) begin
        ds_valid <= 1'b0;
    end
    else if (ds_allowin) begin
        ds_valid <= fs_to_ds_valid;
    end
    /*else if (ws_flush_ds_bus) begin
        ds_valid <= 1'b0;
    end*/
    
    if (fs_to_ds_valid && ds_allowin) begin
        fs_to_ds_bus_r <= fs_to_ds_bus;
    end
end

assign op_31_26  = ds_inst[31:26];
assign op_25_22  = ds_inst[25:22];
assign op_21_20  = ds_inst[21:20];
assign op_19_15  = ds_inst[19:15];

assign rd   = ds_inst[ 4: 0];
assign rj   = ds_inst[ 9: 5];
assign rk   = ds_inst[14:10];

assign i12  = ds_inst[21:10];
assign i20  = ds_inst[24: 5];
assign i16  = ds_inst[25:10];
assign i26  = {ds_inst[ 9: 0], ds_inst[25:10]};

decoder_6_64 u_dec0(.in(op_31_26 ), .out(op_31_26_d ));
decoder_4_16 u_dec1(.in(op_25_22 ), .out(op_25_22_d ));
decoder_2_4  u_dec2(.in(op_21_20 ), .out(op_21_20_d ));
decoder_5_32 u_dec3(.in(op_19_15 ), .out(op_19_15_d ));

assign inst_add_w  = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h00];
assign inst_sub_w  = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h02];
assign inst_slt    = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h04];
assign inst_sltu   = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h05];
assign inst_slti   = op_31_26_d[6'h00] & op_25_22_d[4'h8];
assign inst_sltui  = op_31_26_d[6'h00] & op_25_22_d[4'h9];
assign inst_nor    = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h08];
assign inst_and    = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h09];
assign inst_or     = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h0a];
assign inst_xor    = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h0b];
assign inst_andi   = op_31_26_d[6'h00] & op_25_22_d[4'hd];
assign inst_ori    = op_31_26_d[6'h00] & op_25_22_d[4'he];
assign inst_xori   = op_31_26_d[6'h00] & op_25_22_d[4'hf];
assign inst_slli_w = op_31_26_d[6'h00] & op_25_22_d[4'h1] & op_21_20_d[2'h0] & op_19_15_d[5'h01];
assign inst_srli_w = op_31_26_d[6'h00] & op_25_22_d[4'h1] & op_21_20_d[2'h0] & op_19_15_d[5'h09];
assign inst_srai_w = op_31_26_d[6'h00] & op_25_22_d[4'h1] & op_21_20_d[2'h0] & op_19_15_d[5'h11];
assign inst_sll_w  = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h0e];
assign inst_srl_w  = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h0f];
assign inst_sra_w  = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h10];
assign inst_addi_w = op_31_26_d[6'h00] & op_25_22_d[4'ha];
assign inst_ld_b   = op_31_26_d[6'h0a] & op_25_22_d[4'h0]; 
assign inst_ld_h   = op_31_26_d[6'h0a] & op_25_22_d[4'h1]; 
assign inst_ld_w   = op_31_26_d[6'h0a] & op_25_22_d[4'h2];
assign inst_ld_bu  = op_31_26_d[6'h0a] & op_25_22_d[4'h8];
assign inst_ld_hu  = op_31_26_d[6'h0a] & op_25_22_d[4'h9];
assign inst_st_w   = op_31_26_d[6'h0a] & op_25_22_d[4'h6];
assign inst_st_b   = op_31_26_d[6'h0a] & op_25_22_d[4'h4];
assign inst_st_h   = op_31_26_d[6'h0a] & op_25_22_d[4'h5];
assign inst_jirl   = op_31_26_d[6'h13];
assign inst_b      = op_31_26_d[6'h14];
assign inst_bl     = op_31_26_d[6'h15];
assign inst_beq    = op_31_26_d[6'h16];
assign inst_bne    = op_31_26_d[6'h17];
assign inst_blt    = op_31_26_d[6'h18];
assign inst_bge    = op_31_26_d[6'h19];
assign inst_bltu   = op_31_26_d[6'h1a];
assign inst_bgeu   = op_31_26_d[6'h1b];
assign inst_lu12i_w   = op_31_26_d[6'h05] & ~ds_inst[25];
assign inst_pcaddu12i = op_31_26_d[6'h07] & ~ds_inst[25];
assign inst_mul_w  = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h18];
assign inst_mulh_w = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h19];
assign inst_mulh_wu= op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h1a];
assign inst_div_w  = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h2] & op_19_15_d[5'h00];
assign inst_mod_w  = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h2] & op_19_15_d[5'h01];
assign inst_div_wu = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h2] & op_19_15_d[5'h02];
assign inst_mod_wu = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h2] & op_19_15_d[5'h03];

assign inst_csrrd  = op_31_26_d[6'h01] & ~ds_inst[25] & ~ds_inst[24] & ~|rj;//rj =0
assign inst_csrwr  = op_31_26_d[6'h01] & ~ds_inst[25] & ~ds_inst[24] & (rj == 5'h01);//rj = 1 
assign inst_csrxchg= op_31_26_d[6'h01] & ~ds_inst[25] & ~ds_inst[24] & (rj != 5'h01) & |rj;//rj != 0 & rj != 1
assign inst_ertn   = op_31_26_d[6'h01] & op_25_22_d[4'h9] & op_21_20_d[2'h0] & op_19_15_d[5'h10] & (rk == 5'b01110) & ~|rj & ~|rd;
assign inst_syscall= op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h2] & op_19_15_d[5'h16];
assign inst_break  = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h2] & op_19_15_d[5'h14];
assign inst_rdcntid_w = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h0] & op_19_15_d[5'h00] & (rk == 5'b11000) & ~|rd;
assign inst_rdcntvl_w = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h0] & op_19_15_d[5'h00] & (rk == 5'b11000) & ~|rj;
assign inst_rdcntvh_w = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h0] & op_19_15_d[5'h00] & (rk == 5'b11001) & ~|rj;

//tlb
assign inst_tlbsrch   = op_31_26_d[6'h01] & op_25_22_d[4'h9] & op_21_20_d[2'h0] & op_19_15_d[5'h10] & (rk == 5'b01010) & ~|rj & ~|rd;
assign inst_tlbrd     = op_31_26_d[6'h01] & op_25_22_d[4'h9] & op_21_20_d[2'h0] & op_19_15_d[5'h10] & (rk == 5'b01011) & ~|rj & ~|rd;
assign inst_tlbwr     = op_31_26_d[6'h01] & op_25_22_d[4'h9] & op_21_20_d[2'h0] & op_19_15_d[5'h10] & (rk == 5'b01100) & ~|rj & ~|rd;
assign inst_tlbfill   = op_31_26_d[6'h01] & op_25_22_d[4'h9] & op_21_20_d[2'h0] & op_19_15_d[5'h10] & (rk == 5'b01101) & ~|rj & ~|rd;
assign inst_invtlb    = op_31_26_d[6'h01] & op_25_22_d[4'h9] & op_21_20_d[2'h0] & op_19_15_d[5'h13] & (~|rd[4:3] & ~&rd[2:0]);

assign tlbop = {inst_tlbsrch, inst_tlbrd, inst_tlbwr, inst_tlbfill, inst_invtlb};
assign ex_INE       = ~(inst_add_w | inst_sub_w | inst_addi_w |
                        inst_slt | inst_sltu | inst_slti | inst_sltui | 
                        inst_nor | inst_and | inst_or | inst_xor | inst_andi |inst_ori | inst_xori | 
                        inst_sll_w | inst_srl_w | inst_sra_w | inst_slli_w | inst_srli_w | inst_srai_w|
                        inst_ld_b | inst_ld_h | inst_ld_w | inst_ld_bu | inst_ld_hu |
                        inst_st_b | inst_st_h | inst_st_w|
                        inst_jirl | inst_b | inst_bl | inst_beq | inst_bne | inst_blt | inst_bge | inst_bltu | inst_bgeu |
                        inst_lu12i_w | inst_pcaddu12i |
                        inst_mul_w | inst_mulh_w | inst_mulh_wu |
                        inst_div_w | inst_div_wu | inst_mod_w | inst_mod_wu |
                        inst_csrrd | inst_csrwr | inst_csrxchg | inst_ertn | inst_syscall | inst_break |
                        inst_rdcntid_w | inst_rdcntvl_w | inst_rdcntvh_w |
                        inst_tlbsrch | inst_tlbrd   | inst_tlbwr  | inst_tlbfill   | (inst_invtlb && invtlb_op<7)
                        );
assign csr_we       = inst_csrwr | inst_csrxchg;
assign csr_re       = inst_csrwr | inst_csrrd | inst_csrxchg | inst_rdcntid_w;
assign csr_wmask    = inst_csrxchg ? rj_value : {32{1'b1}};
assign csr_num      = inst_rdcntid_w ? `CSR_TID : ds_inst[23:10];
assign inst_cnt_op  = {3{inst_rdcntid_w}} & 3'b001 |
                      {3{inst_rdcntvl_w}} & 3'b010 |
                      {3{inst_rdcntvh_w}} & 3'b100 ;
assign inst_st_op = {3{inst_st_b}} & 3'b001
                   |{3{inst_st_h}} & 3'b010
                   |{3{inst_st_w}} & 3'b100;
                   
assign inst_ld_op = {5{inst_ld_b}} & 5'b00001
                   |{5{inst_ld_h}} & 5'b00010
                   |{5{inst_ld_w}} & 5'b00100
                   |{5{inst_ld_bu}}& 5'b01000
                   |{5{inst_ld_hu}}& 5'b10000;

assign invtlb_op = ds_inst[4:0];        
          
assign alu_op[ 0] = inst_add_w | inst_addi_w | inst_ld_w | inst_ld_b | inst_ld_h
                    |inst_ld_bu | inst_ld_hu | inst_st_w | inst_st_b | inst_st_h
                    | inst_jirl | inst_bl | inst_pcaddu12i;
assign alu_op[ 1] = inst_sub_w;
assign alu_op[ 2] = inst_slt  | inst_slti;
assign alu_op[ 3] = inst_sltu | inst_sltui;
assign alu_op[ 4] = inst_and  | inst_andi;
assign alu_op[ 5] = inst_nor;
assign alu_op[ 6] = inst_or   | inst_ori;
assign alu_op[ 7] = inst_xor  | inst_xori;
assign alu_op[ 8] = inst_slli_w | inst_sll_w;
assign alu_op[ 9] = inst_srli_w | inst_srl_w;
assign alu_op[10] = inst_srai_w | inst_sra_w;
assign alu_op[11] = inst_lu12i_w;
assign alu_op[12] = inst_mul_w;
assign alu_op[13] = inst_mulh_w;
assign alu_op[14] = inst_mulh_wu;
assign alu_op[15] = inst_div_w;
assign alu_op[16] = inst_mod_w;
assign alu_op[17] = inst_div_wu;
assign alu_op[18] = inst_mod_wu;

assign need_ui5   =  inst_slli_w | inst_srli_w | inst_srai_w;
assign need_si12  =  inst_addi_w | inst_ld_w | inst_ld_b | inst_ld_h | inst_ld_bu
                    | inst_ld_hu | inst_st_w | inst_st_b | inst_st_h | inst_slti | inst_sltui;
assign need_ui12  =  inst_andi | inst_ori | inst_xori;
assign need_si16  =  inst_jirl | inst_beq | inst_bne | inst_blt 
                    | inst_bge | inst_bltu | inst_bgeu;
assign need_si20  =  inst_lu12i_w | inst_pcaddu12i;
assign need_si26  =  inst_b | inst_bl;
assign src2_is_4  =  inst_jirl | inst_bl;


assign ds_imm = src2_is_4 ? 32'h4                      :
		        need_si20 ? {i20[19:0], 12'b0}         :  //i20[16:5]==i12[11:0]
                need_ui12 ? {20'b0, i12[11:0]}         :
                            {{20{i12[11]}}, i12[11:0]} ;  /*need_ui5 || need_si12*/

assign br_offs = need_si26 ? {{ 4{i26[25]}}, i26[25:0], 2'b0} : 
                             {{14{i16[15]}}, i16[15:0], 2'b0} ;

assign jirl_offs = {{14{i16[15]}}, i16[15:0], 2'b0};

assign src_reg_is_rd = inst_beq | inst_bne | inst_blt | inst_bge | inst_bltu | inst_bgeu 
                    | inst_st_w | inst_st_b| inst_st_h|inst_csrwr| inst_csrxchg;

assign src1_is_pc    = inst_jirl | inst_bl | inst_pcaddu12i;

assign src2_is_imm   = inst_slli_w | 
                       inst_srli_w |
                       inst_srai_w |
                       inst_addi_w |
                       inst_ld_w   |
                       inst_ld_b   |
                       inst_ld_h   |
                       inst_ld_bu  |
                       inst_ld_hu  |
                       inst_st_w   |
                       inst_st_b   |
                       inst_st_h   |
                       inst_lu12i_w|
                       inst_jirl   |
                       inst_bl     |
                       inst_slti   |
                       inst_sltui  |
                       inst_andi   |
                       inst_ori    |
                       inst_xori   |
                       inst_pcaddu12i;


assign res_from_mem  = inst_ld_w | inst_ld_b | inst_ld_h | inst_ld_bu | inst_ld_hu;
assign dst_is_r1     = inst_bl;
assign gr_we         = ~inst_st_w & ~inst_beq & ~inst_bne & ~inst_b & ~inst_st_b
                        & ~inst_st_h & ~inst_blt & ~inst_bge & ~inst_bltu & ~inst_bgeu
                        & ~inst_ertn & ~inst_syscall & ~inst_break & ~ex_INE 
                        & ~inst_tlbsrch & ~inst_tlbrd & ~inst_tlbwr & ~inst_tlbfill &~inst_invtlb;
assign mem_we        = inst_st_w | inst_st_b |inst_st_h;
assign dest          = dst_is_r1 ? 5'd1 :
                       inst_rdcntid_w ? rj : rd;


assign raddr1_valid = (inst_add_w |   // inst
                       inst_sub_w |
                       inst_addi_w|
                       inst_beq   |
                       inst_bne   |
                       inst_blt   |
                       inst_bge   |
                       inst_bltu  |
                       inst_bgeu  |
                       inst_jirl  |
                       inst_slt   |
                       inst_sltu  |
                       inst_slti  |
                       inst_sltui |
                       inst_and   |
                       inst_or    |
                       inst_xor   |
                       inst_nor   |
                       inst_andi  |
                       inst_ori   |
                       inst_xori  |
                       inst_sll_w |
                       inst_srl_w |
                       inst_sra_w |
                       inst_slli_w|
                       inst_srli_w|
                       inst_srai_w|
                       inst_ld_w  |
                       inst_ld_b  |
                       inst_ld_h  |
                       inst_ld_bu |
                       inst_ld_hu |
                       inst_st_w  |
                       inst_st_b  |
                       inst_st_h  |
                       inst_mul_w |
                       inst_mulh_w|
                       inst_mulh_wu|
                       inst_div_w  |
                       inst_mod_w  |
                       inst_div_wu |
                       inst_mod_wu |
                       inst_csrxchg|
                       inst_invtlb
                      ) & (|rf_raddr1) // rf_raddr1 != 0
                        & ds_valid; 

assign raddr2_valid = (inst_add_w |   // inst
                       inst_sub_w |
                       inst_beq   |
                       inst_bne   |
                       inst_blt   |
                       inst_bge   |
                       inst_bltu  |
                       inst_bgeu  |
                       inst_slt   |
                       inst_sltu  |
                       inst_and   |
                       inst_or    |
                       inst_xor   |
                       inst_nor   |
                       inst_sll_w |
                       inst_srl_w |
                       inst_sra_w |
                       inst_st_w  |
                       inst_st_b  |
                       inst_st_h  |
                       inst_mul_w |
                       inst_mulh_w|
                       inst_mulh_wu|
                       inst_div_w  |
                       inst_mod_w  |
                       inst_div_wu |
                       inst_mod_wu |
                       inst_csrwr  |
                       inst_csrxchg|
                       inst_invtlb 
                      ) & (|rf_raddr2) // rf_raddr1 != 0
                        & ds_valid; 


assign rf_raddr1 = rj;
assign rf_raddr2 = src_reg_is_rd ? rd :rk;
regfile u_regfile(
    .clk    (clk      ),
    .raddr1 (rf_raddr1),
    .rdata1 (rf_rdata1),
    .raddr2 (rf_raddr2),
    .rdata2 (rf_rdata2),
    .we     (rf_we    ),
    .waddr  (rf_waddr ),
    .wdata  (rf_wdata )
    );

assign es_read1_unuse   =  es_relate_r1 && es_read_except;
assign es_read2_unuse   =  es_relate_r2 && es_read_except;
assign ms_read1_unuse   =  ms_relate_r1 && ms_read_except;
assign ms_read2_unuse   =  ms_relate_r2 && ms_read_except;
assign ds_ready_go = ~(es_read1_unuse | es_read2_unuse | ms_read1_unuse | ms_read2_unuse);

assign es_relate_r1 = (rf_raddr1 == es_dest) && es_dest_valid && raddr1_valid;
assign es_relate_r2 = (rf_raddr2 == es_dest) && es_dest_valid && raddr2_valid;
assign ms_relate_r1 = (rf_raddr1 == ms_dest) && ms_dest_valid && raddr1_valid;
assign ms_relate_r2 = (rf_raddr2 == ms_dest) && ms_dest_valid && raddr2_valid;
assign ws_relate_r1 = (rf_raddr1 == ws_dest) && ws_dest_valid && raddr1_valid;
assign ws_relate_r2 = (rf_raddr2 == ws_dest) && ws_dest_valid && raddr2_valid;

assign rj_value  =   es_relate_r1 ? es_to_ds_bus :
                    (ms_relate_r1 ? ms_to_ds_bus :
                    (ws_relate_r1 ? ws_to_ds_bus :
                     rf_rdata1));

assign rkd_value =   es_relate_r2 ? es_to_ds_bus :
                    (ms_relate_r2 ? ms_to_ds_bus :
                    (ws_relate_r2 ? ws_to_ds_bus :
                     rf_rdata2));

assign rj_eq_rd = rj_value == rkd_value;
assign rj_le_rd = $signed(rj_value) < $signed(rkd_value);
assign rj_leu_rd = rj_value < rkd_value;

assign br_inst_valid = (   inst_beq  &&  rj_eq_rd
                   || inst_bne  && !rj_eq_rd
                   || inst_blt  &&  rj_le_rd
                   || inst_bge  && !rj_le_rd
                   || inst_bltu &&  rj_leu_rd
                   || inst_bgeu && !rj_leu_rd
                   || inst_jirl
                   || inst_bl
                   || inst_b
                  ) && ds_valid;
assign br_stall = br_inst_valid && es_inst_load && (es_relate_r1 || es_relate_r2);
assign br_taken = br_inst_valid && ds_ready_go ;//&& !ws_flush_ds_bus; 
assign br_target = (inst_beq || inst_bne || inst_blt || inst_bge || inst_bltu 
                 || inst_bgeu|| inst_bl || inst_b) ? (ds_pc + br_offs) :
                                     /*inst_jirl*/ (rj_value + jirl_offs);

endmodule